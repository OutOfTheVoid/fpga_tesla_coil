module GateDrivePhaser (
	input 
);